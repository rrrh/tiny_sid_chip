VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO svf_2nd
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN svf_2nd 0 0 ;
  SIZE 62.000 BY 72.000 ;
  SYMMETRY X Y ;

  PIN vin
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 34.000 0.500 38.000 ;
    END
  END vin

  PIN vout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 61.500 34.000 62.000 38.000 ;
    END
  END vout

  PIN sel0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 9.000 0.500 11.000 ;
    END
  END sel0

  PIN sel1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 15.000 0.500 17.000 ;
    END
  END sel1

  PIN sc_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 51.000 0.500 53.000 ;
    END
  END sc_clk

  PIN q0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 55.000 0.500 57.000 ;
    END
  END q0

  PIN q1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 57.000 0.500 59.000 ;
    END
  END q1

  PIN q2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 59.000 0.500 61.000 ;
    END
  END q2

  PIN q3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 61.000 0.500 63.000 ;
    END
  END q3

  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 70.000 62.000 72.000 ;
    END
  END vdd

  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 0.000 62.000 2.000 ;
    END
  END vss

  OBS
    LAYER Metal1 ;
      RECT 0.500 0.500 61.500 71.500 ;
    LAYER Metal2 ;
      RECT 0.500 0.500 61.500 71.500 ;
  END

END svf_2nd

END LIBRARY
