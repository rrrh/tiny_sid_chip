VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO r2r_dac_8bit
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN r2r_dac_8bit 0 0 ;
  SIZE 38.000 BY 45.000 ;
  SYMMETRY X Y ;

  PIN d0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 2.500 0.500 3.500 ;
    END
  END d0

  PIN d1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 6.500 0.500 7.500 ;
    END
  END d1

  PIN d2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 10.500 0.500 11.500 ;
    END
  END d2

  PIN d3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 14.500 0.500 15.500 ;
    END
  END d3

  PIN d4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 18.500 0.500 19.500 ;
    END
  END d4

  PIN d5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 22.500 0.500 23.500 ;
    END
  END d5

  PIN d6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 26.500 0.500 27.500 ;
    END
  END d6

  PIN d7
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 30.500 0.500 31.500 ;
    END
  END d7

  PIN vout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 37.500 20.500 38.000 21.500 ;
    END
  END vout

  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 43.000 38.000 45.000 ;
    END
  END vdd

  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 0.000 38.000 2.000 ;
    END
  END vss

  OBS
    LAYER Metal1 ;
      RECT 0.500 0.500 37.500 44.500 ;
    LAYER Metal2 ;
      RECT 0.500 0.500 37.500 44.500 ;
  END

END r2r_dac_8bit

END LIBRARY
