VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO svf_2nd
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN svf_2nd 0 0 ;
  SIZE 62.000 BY 68.000 ;
  SYMMETRY X Y ;

  PIN vin
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 32.000 0.500 36.000 ;
    END
  END vin

  PIN vout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 61.500 32.000 62.000 36.000 ;
    END
  END vout

  PIN sel0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 9.000 0.500 11.000 ;
    END
  END sel0

  PIN sel1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 15.000 0.500 17.000 ;
    END
  END sel1

  PIN sc_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 48.000 0.500 50.000 ;
    END
  END sc_clk

  PIN q0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 52.000 0.500 54.000 ;
    END
  END q0

  PIN q1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 54.000 0.500 56.000 ;
    END
  END q1

  PIN q2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 56.000 0.500 58.000 ;
    END
  END q2

  PIN q3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 58.000 0.500 60.000 ;
    END
  END q3

  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 66.000 62.000 68.000 ;
    END
  END vdd

  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 0.000 62.000 2.000 ;
    END
  END vss

  OBS
    LAYER Metal1 ;
      RECT 0.500 0.500 61.500 67.500 ;
    LAYER Metal2 ;
      RECT 0.500 0.500 61.500 67.500 ;
  END

END svf_2nd

END LIBRARY
