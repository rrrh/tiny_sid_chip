VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sar_adc_8bit
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sar_adc_8bit 0 0 ;
  SIZE 42.000 BY 45.000 ;
  SYMMETRY X Y ;

  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 4.500 0.500 5.500 ;
    END
  END clk

  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 8.500 0.500 9.500 ;
    END
  END rst_n

  PIN vin
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 21.500 0.500 22.500 ;
    END
  END vin

  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 12.500 0.500 13.500 ;
    END
  END start

  PIN eoc
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 41.500 4.500 42.000 5.500 ;
    END
  END eoc

  PIN dout0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 41.500 8.500 42.000 9.500 ;
    END
  END dout0

  PIN dout1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 41.500 13.000 42.000 14.000 ;
    END
  END dout1

  PIN dout2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 41.500 17.500 42.000 18.500 ;
    END
  END dout2

  PIN dout3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 41.500 22.000 42.000 23.000 ;
    END
  END dout3

  PIN dout4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 41.500 26.500 42.000 27.500 ;
    END
  END dout4

  PIN dout5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 41.500 31.000 42.000 32.000 ;
    END
  END dout5

  PIN dout6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 41.500 35.500 42.000 36.500 ;
    END
  END dout6

  PIN dout7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 41.500 40.000 42.000 41.000 ;
    END
  END dout7

  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 43.000 42.000 45.000 ;
    END
  END vdd

  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 0.000 42.000 2.000 ;
    END
  END vss

  OBS
    LAYER Metal1 ;
      RECT 0.500 0.500 41.500 44.500 ;
    LAYER Metal2 ;
      RECT 0.500 0.500 41.500 44.500 ;
  END

END sar_adc_8bit

END LIBRARY
