VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO r2r_dac_8bit
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN r2r_dac_8bit 0 0 ;
  SIZE 38.000 BY 48.000 ;
  SYMMETRY X Y ;

  PIN d0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3.000 0.500 4.000 ;
    END
  END d0

  PIN d1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 8.000 0.500 9.000 ;
    END
  END d1

  PIN d2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 13.000 0.500 14.000 ;
    END
  END d2

  PIN d3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 18.000 0.500 19.000 ;
    END
  END d3

  PIN d4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 23.000 0.500 24.000 ;
    END
  END d4

  PIN d5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 28.000 0.500 29.000 ;
    END
  END d5

  PIN d6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 33.000 0.500 34.000 ;
    END
  END d6

  PIN d7
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 38.000 0.500 39.000 ;
    END
  END d7

  PIN vout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 37.500 23.500 38.000 24.500 ;
    END
  END vout

  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 46.000 38.000 48.000 ;
    END
  END vdd

  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 0.000 38.000 2.000 ;
    END
  END vss

  OBS
    LAYER Metal1 ;
      RECT 0.500 0.500 37.500 47.500 ;
    LAYER Metal2 ;
      RECT 0.500 0.500 37.500 47.500 ;
  END

END r2r_dac_8bit

END LIBRARY
