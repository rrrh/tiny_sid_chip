VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO bias_dac_2ch
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN bias_dac_2ch 0 0 ;
  SIZE 35.000 BY 40.000 ;
  SYMMETRY X Y ;

  PIN dfc0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 23.500 0.500 24.500 ;
    END
  END dfc0

  PIN dfc1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 27.000 0.500 28.000 ;
    END
  END dfc1

  PIN dfc2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 30.500 0.500 31.500 ;
    END
  END dfc2

  PIN dfc3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 34.000 0.500 35.000 ;
    END
  END dfc3

  PIN dq0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 3.500 0.500 4.500 ;
    END
  END dq0

  PIN dq1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 7.000 0.500 8.000 ;
    END
  END dq1

  PIN dq2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 10.500 0.500 11.500 ;
    END
  END dq2

  PIN dq3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 14.000 0.500 15.000 ;
    END
  END dq3

  PIN vout_fc
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 34.500 29.500 35.000 30.500 ;
    END
  END vout_fc

  PIN vout_q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 34.500 11.500 35.000 12.500 ;
    END
  END vout_q

  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 38.000 35.000 40.000 ;
    END
  END vdd

  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 0.000 35.000 2.000 ;
    END
  END vss

  OBS
    LAYER Metal1 ;
      RECT 0.500 0.500 34.500 39.500 ;
    LAYER Metal2 ;
      RECT 0.500 0.500 34.500 39.500 ;
  END

END bias_dac_2ch

END LIBRARY
