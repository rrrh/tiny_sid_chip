VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sar_adc_8bit
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sar_adc_8bit 0 0 ;
  SIZE 42.000 BY 42.000 ;
  SYMMETRY X Y ;

  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 4.500 0.500 5.500 ;
    END
  END clk

  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 8.500 0.500 9.500 ;
    END
  END rst_n

  PIN vin
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 19.500 0.500 20.500 ;
    END
  END vin

  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 12.500 0.500 13.500 ;
    END
  END start

  PIN eoc
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 41.500 4.500 42.000 5.500 ;
    END
  END eoc

  PIN dout0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 41.500 7.500 42.000 8.500 ;
    END
  END dout0

  PIN dout1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 41.500 11.000 42.000 12.000 ;
    END
  END dout1

  PIN dout2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 41.500 14.500 42.000 15.500 ;
    END
  END dout2

  PIN dout3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 41.500 18.000 42.000 19.000 ;
    END
  END dout3

  PIN dout4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 41.500 21.500 42.000 22.500 ;
    END
  END dout4

  PIN dout5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 41.500 25.000 42.000 26.000 ;
    END
  END dout5

  PIN dout6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 41.500 28.500 42.000 29.500 ;
    END
  END dout6

  PIN dout7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 41.500 32.000 42.000 33.000 ;
    END
  END dout7

  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 40.000 42.000 42.000 ;
    END
  END vdd

  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 0.000 42.000 2.000 ;
    END
  END vss

  OBS
    LAYER Metal1 ;
      RECT 0.500 0.500 41.500 41.500 ;
    LAYER Metal2 ;
      RECT 0.500 0.500 41.500 41.500 ;
  END

END sar_adc_8bit

END LIBRARY
