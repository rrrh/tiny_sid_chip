VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sar_adc_8bit
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sar_adc_8bit 0 0 ;
  SIZE 95.000 BY 104.000 ;
  SYMMETRY X Y ;

  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 8.000 0.500 9.000 ;
    END
  END clk

  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 14.000 0.500 15.000 ;
    END
  END rst_n

  PIN vin
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 52.000 0.500 53.000 ;
    END
  END vin

  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 20.000 0.500 21.000 ;
    END
  END start

  PIN eoc
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.500 8.000 95.000 9.000 ;
    END
  END eoc

  PIN dout[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.500 18.000 95.000 19.000 ;
    END
  END dout[0]

  PIN dout[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.500 24.000 95.000 25.000 ;
    END
  END dout[1]

  PIN dout[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.500 30.000 95.000 31.000 ;
    END
  END dout[2]

  PIN dout[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.500 36.000 95.000 37.000 ;
    END
  END dout[3]

  PIN dout[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.500 42.000 95.000 43.000 ;
    END
  END dout[4]

  PIN dout[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.500 48.000 95.000 49.000 ;
    END
  END dout[5]

  PIN dout[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.500 54.000 95.000 55.000 ;
    END
  END dout[6]

  PIN dout[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.500 60.000 95.000 61.000 ;
    END
  END dout[7]

  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 102.000 95.000 104.000 ;
    END
  END vdd

  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 0.000 95.000 2.000 ;
    END
  END vss

  OBS
    LAYER Metal1 ;
      RECT 0.500 0.500 94.500 103.500 ;
    LAYER Metal2 ;
      RECT 0.500 0.500 94.500 103.500 ;
  END

END sar_adc_8bit

END LIBRARY
